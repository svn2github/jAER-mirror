package settings is
	constant FX3_CLOCK_FREQ : integer := 100;
	constant FX3_EARLY_PACKET_MS : integer := 1;
	constant LOGIC_CLOCK_FREQ : integer := 25;
end settings;

