library ieee;
use ieee.std_logic_1164.all;

entity ExtTriggerSPIConfig is
	port (
		Clock_CI : in std_logic;
		Reset_RI : in std_logic);
end entity ExtTriggerSPIConfig;

architecture Behavioral of ExtTriggerSPIConfig is
	
begin

end architecture Behavioral;
