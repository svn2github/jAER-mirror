library ieee;
use ieee.std_logic_1164.all;

entity APSADCSPIConfig is
	port (
		Clock_CI : in std_logic;
		Reset_RI : in std_logic);
end entity APSADCSPIConfig;

architecture Behavioral of APSADCSPIConfig is
	
begin

end architecture Behavioral;
