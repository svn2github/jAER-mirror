--------------------------------------------------------------------------------
-- Company: INI
-- Engineer: Diederik Paul Moeys
--
-- Create Date:    28.08.2014
-- Design Name:    
-- Module Name:    MullerCelement
-- Project Name:   VISUALISE
-- Target Device:  Latticed LFE3-17EA-7ftn256i
-- Tool versions:  Diamond x64 3.0.0.97x
-- Description:	   Mueller C-element
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Libraries -------------------------------------------------------------------
-------------------------------------------------------------------------------- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Entity Declaration ----------------------------------------------------------
--------------------------------------------------------------------------------
entity MullerCelement is
	port (
	Ain,Bin : 	in	std_logic; 
	Cout 	: 	out std_logic);
end MullerCelement;
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Architecture Declaration ----------------------------------------------------
--------------------------------------------------------------------------------
architecture Behavioural of MullerCelement is
begin
process (Ain, Bin)
    variable state  : std_logic;
    variable in_cat : std_logic_vector (1 downto 0);
begin
	in_cat := (Ain, Bin);
	case (in_cat) is
		when "00" =>  state := '0';
		when "01" =>  state := state;
		when "10" =>  state := state;
		when "11" =>  state := '1';
		when others => null;
    end case;
	Cout <= state;
end process;
end Behavioural;
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------