library ieee;
use ieee.std_logic_1164.all;

entity BiasGenStateMachine is
	port (
		Clock_CI : in std_logic;
		Reset_RI : in std_logic
	);
end entity BiasGenStateMachine;

architecture Behavioral of BiasGenStateMachine is
	
begin
	
end architecture Behavioral;
